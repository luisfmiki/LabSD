LIBRARY IEEE;
use ieee.std_logic_1164.all;

entity FlipFlopD is
	port( clk: in std_logic;
		  D: in std_logic;
	      Q: out std_logic;
			reset: in std_logic
	    );
end FlipFlopD;

architecture RTL of FlipFlopD is
begin
	Q <= 
	'0' when (reset='1') else
	D when rising_edge(clk);
	
	
--	process(clock)
--	begin
--		if (clock='1' and clock'event) then
--			Q <= D;
--		end if;
--	end process;
end RTL;

