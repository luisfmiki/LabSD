LIBRARY IEEE;
use ieee.std_logic_1164.all;

entity tb_Mux is
end tb_Mux;
architecture teste of tb_Mux is
component Mux is
port ( A,R,S: in std_logic;
F: out std_logic);

end component;

	signal fio_A, fio_R: std_logic;
	signal fio_S, fio_F: std_logic;
begin
instancia_Mux: Mux port map(A=>fio_A, R=>fio_R, S=>fio_S,
F=>fio_F);
fio_A <= '1' after 5ns; 
fio_R <= '0' after 5ns;
fio_S <= '0' after 3ns, '1' after 7ns;

end teste;